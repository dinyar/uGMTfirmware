-- ipbus_dpram_asym
--
-- Generic dual-port memory with asymmetric port widths and ipbus access on one
-- port. Requires data file with one value per line in hexadecimal notation (no
-- '0x' though) for initialization.
--
-- Should lead to an inferred block RAM in Xilinx parts with modern tools
--
-- Note the wait state on ipbus access - full speed access is not possible
-- Can combine with peephole_ram access method for full speed access.
--
-- Dave Newbold, July 2013
-- Dinyar Rabady, March 2015

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use work.ipbus.all;

use STD.TEXTIO.all;
use ieee.std_logic_textio.all;

entity ipbus_dpram_asym is
	generic(
		DATA_FILE: string;
		ADDR_WIDTH: natural;
		WORD_WIDTH: natural := 32
	);
	port(
		clk: in std_logic;
		rst: in std_logic;
		ipb_in: in ipb_wbus;
		ipb_out: out ipb_rbus;
		rclk: in std_logic;
		we: in std_logic := '0';
		d: in std_logic_vector(31 downto 0) := (others => '0');
		q: out std_logic_vector(WORD_WIDTH - 1 downto 0);
		addr: in std_logic_vector(ADDR_WIDTH - 1 downto 0)
	);

end ipbus_dpram_asym;

architecture rtl of ipbus_dpram_asym is

	-- TODO: Is there a less stupid way to compute those two values?
	-- (i.e.: can I write one function that does this?)
	function find_ipbus_addr_width (algo_word_width : integer; algo_addr_width : integer) return natural is
		variable ipb_word_width : natural := algo_word_width;
		variable ipb_addr_width : natural := algo_addr_width;
	begin
		-- If word size is 16 it will be doubled to 32 in the last iteration.
		while ipb_word_width <= 16 loop
			ipb_word_width := ipb_word_width * 2;
			ipb_addr_width := ipb_addr_width - 1;
		end loop;
		return ipb_addr_width;
	end function find_ipbus_addr_width;
	function find_ipbus_word_width (algo_word_width : integer; algo_addr_width : integer) return natural is
		variable ipb_word_width : natural := algo_word_width;
		variable ipb_addr_width : natural := algo_addr_width;
	begin
		-- If word size is 16 it will be doubled to 32 in the last iteration.
		while ipb_word_width <= 16 loop
			ipb_word_width := ipb_word_width * 2;
			ipb_addr_width := ipb_addr_width - 1;
		end loop;
		return ipb_word_width;
	end function find_ipbus_word_width;

	constant ALGO_WORD_SIZE : natural := WORD_WIDTH;
	constant ALGO_ADDR_WIDTH : natural := ADDR_WIDTH;
	constant IPBUS_WORD_SIZE : natural := find_ipbus_word_width(ALGO_WORD_SIZE, ALGO_ADDR_WIDTH);
	constant IPBUS_ADDR_WIDTH : natural := find_ipbus_addr_width(ALGO_WORD_SIZE, ALGO_ADDR_WIDTH);
	constant ratio : integer := IPBUS_WORD_SIZE/ALGO_WORD_SIZE;

	function log2 (val : integer) return natural is
		variable res : natural;
	begin
		for i in 0 to 31 loop
			if (val <= (2**i)) then
				res := i;
				exit;
			end if;
		end loop;
		return res;
	end function log2;


	-- Direction of array important to make first word in data file correspond
	-- to first address.
	type ram_array is array(0 to 2 ** ALGO_ADDR_WIDTH - 1) of std_logic_vector(ALGO_WORD_SIZE - 1 downto 0);

    impure function InitRamFromFile (file_name : in string) return ram_array is
        file F : text open read_mode is file_name;
        variable L : line;
        variable ram : ram_array;
    begin
        for i in ram_array'range loop
            readline (F, L);
            hread (L, ram(i));
        end loop;
        return ram;
    end function;

	shared variable ram: ram_array := InitRamFromFile(DATA_FILE);

	signal sel : integer range 0 to 2 ** IPBUS_ADDR_WIDTH - 1 := 0;
	signal rsel: integer range 0 to 2 ** ALGO_ADDR_WIDTH - 1 := 0;
	signal ack: std_logic;

    signal reduced_ipbus_in, reduced_ipbus_out : std_logic_vector(IPBUS_WORD_SIZE - 1 downto 0);

begin

	sel <= to_integer(unsigned(ipb_in.ipb_addr(IPBUS_ADDR_WIDTH - 1 downto 0)));
	reduced_ipbus_in <= ipb_in.ipb_wdata(IPBUS_WORD_SIZE - 1 downto 0);

	process(clk)
	begin
		if rising_edge(clk) then
			for i in 0 to ratio - 1 loop

				reduced_ipbus_out((i+1)*ALGO_WORD_SIZE - 1 downto i*ALGO_WORD_SIZE)
					<= ram(to_integer(
						unsigned(ipb_in.ipb_addr(IPBUS_ADDR_WIDTH - 1 downto 0)) & to_unsigned(i, log2(ratio))
				)); -- Order of statements is important to infer read-first RAM!

				if ipb_in.ipb_strobe='1' and ipb_in.ipb_write='1' then

					ram(to_integer(
						unsigned(ipb_in.ipb_addr(IPBUS_ADDR_WIDTH - 1 downto 0)) & to_unsigned(i, log2(ratio))
					)) := reduced_ipbus_in( (i+1)*ALGO_WORD_SIZE - 1 downto i*ALGO_WORD_SIZE );

				end if;
			end loop;
			ack <= ipb_in.ipb_strobe and not ack;
		end if;
	end process;

	ipb_out.ipb_rdata(IPBUS_WORD_SIZE - 1 downto 0) <= reduced_ipbus_out;
	ipb_out.ipb_ack <= ack;
	ipb_out.ipb_err <= '0';

	rsel <= to_integer(unsigned(addr));

	process(rclk)
	begin
		if rising_edge(rclk) then
			q <= ram(rsel); -- Order of statements is important to infer read-first RAM!
			if we = '1' then
				ram(rsel) := d;
			end if;
		end if;
	end process;

end rtl;
